`timescale 1ns/1ps
`include "./sub_64bit.v"
`include "../ADD/add_64bit.v"

module sub_64bit_tb;

    reg signed [63:0] a;
    reg signed [63:0] b;
    wire signed [63:0] out;
    wire overflow;

    sub_64bit f1(a, b, out, overflow);

    initial begin
        $dumpfile("sub_64bit_tb.vcd");
        $dumpvars(0, sub_64bit_tb);

        $monitor("a\t= %b\t%d\nb\t= %b\t%d\nout\t= %b\t%d\noverflow= %d\n", a, a, b, b, out, out, overflow);

        b = 64'b1000000000000000000000000000000000000000000000000000000000000000;
        a = 64'b1111111111111111111111111111111111111111111111111111111111111111;

        a = 64'b0111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111;
        b = 64'b0111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111;

        #10
        a = 64'b1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
        b = 64'b1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;

        #10
        a = 64'b0111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111;
        b = 64'b1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;

        #10
        a = 64'b1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
        b = 64'b0111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111;

        #10
        a = 64'b0101;
        b = 64'b1110;

    end

endmodule