`timescale 1ns/1ps
`include "alu.v"

module alu_tb;

    reg signed [63:0] a;
    reg signed [63:0] b;
    wire signed [63:0] out;
    wire overflow;
    reg [1:0] control;

    alu f(control, a, b, out, overflow);

    initial begin
        $dumpfile("alu_tb.vcd");
        $dumpvars(0, alu_tb);

        a=64'b0000000000000000000000000000000000000000000000000000000000000000;
		b=64'b0000000000000000000000000000000000000000000000000000000000000000;

		control = 2'b11;

        $monitor("Control = %d\na   = %b\t%d\nb   = %b\t%d\nout = %b\t%d\nOverflow = %d\n", control, a, a, b, b, out, out, overflow);

        #10
        a = 64'b0111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111;
        b = 64'b0111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111;

        #10
        a = 64'b1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
        b = 64'b1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;

        #10
        a = 64'b0111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111;
        b = 64'b1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;

        #10
        a = 64'b1000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
        b = 64'b0111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111_1111;
    end

endmodule